library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;

-- entidade do testbench
entity random_generator_tb is
end entity;

architecture tb of random_generator_tb is
     